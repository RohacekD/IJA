�� sr ija.ija2015.homework2.game.Game��T��}"� Z endedZ otherCantPlayL blackPlayert #Lija/ija2015/homework2/game/Player;L boardt #Lija/ija2015/homework2/board/Board;[ countst [IL currentPlayerq ~ L whitePlayerq ~ xp  sr #ija.ija2015.homework2.game.AiPlayerހ�>{�wQ L aiTypet &Lija/ija2015/homework2/game/Player$Ai;xr !ija.ija2015.homework2.game.Player�^품zU� Z alreadyCheckedI countOfDiskZ initializedI takenFromPoolZ whiteL legalst Ljava/util/ArrayList;[ poolt #[Lija/ija2015/homework2/board/Disk;L 
toTurnOverq ~ xp       sr java.util.ArrayListx����a� I sizexp   w   sr &ija.ija2015.homework2.board.BoardField�7*����� I colsI rowL diskt "Lija/ija2015/homework2/board/Disk;[ surroundingt $[Lija/ija2015/homework2/board/Field;xp      pur $[Lija.ija2015.homework2.board.Field;'m' 0VA  xp   sq ~       sr  ija.ija2015.homework2.board.DiskJ�~j��U~ Z isWhitexpuq ~    sr 'ija.ija2015.homework2.board.BorderField��C̈��  xpsq ~ sq ~ sq ~       sq ~ uq ~    q ~ q ~ sq ~ sq ~ sq ~ q ~ sq ~       sq ~ uq ~    sq ~       sq ~ uq ~    sq ~ q ~ q ~ q ~ q ~ !sq ~       sq ~  uq ~    sq ~ q ~ $q ~ q ~ !sq ~       puq ~    q ~ (q ~ !q ~ sq ~       puq ~    q ~ !q ~ q ~  sq ~ sq ~ sq ~ sq ~ q ~ ,q ~ 2q ~ 3sq ~ sq ~       puq ~    sq ~ q ~ (q ~ !q ~ ,q ~ 3q ~ 4sq ~ sq ~ q ~ 5q ~ 9q ~ 7q ~ 7q ~ +q ~ q ~ q ~ q ~ .q ~ ,q ~ 5q ~ (q ~ q ~ q ~ !q ~ (q ~ $q ~ q ~ q ~  q ~ 0q ~ .q ~ ,q ~ !xur #[Lija.ija2015.homework2.board.Disk;���ɦ��  xp   q ~ q ~ )sq ~  sq ~  sq ~     w    x~r $ija.ija2015.homework2.game.Player$Ai          xr java.lang.Enum          xpt humansr !ija.ija2015.homework2.board.Boardzg`8��j [ deskt %[[Lija/ija2015/homework2/board/Field;L rulest #Lija/ija2015/homework2/board/Rules;xpur %[[Lija.ija2015.homework2.board.Field;�z��T(�  xp   uq ~    q ~ 'q ~ q ~ q ~ q ~ uq ~    q ~ +q ~ $q ~ q ~ q ~ uq ~    q ~ 7q ~ (q ~ !q ~ q ~  uq ~    q ~ 9q ~ 5q ~ ,q ~ .q ~ 0uq ~    q ~ 8q ~ 4q ~ 3q ~ 2q ~ 1sr 'ija.ija2015.homework2.game.ReversiRuless��7ŗ/ I sizexp   ur [IM�`&v겥  xp         q ~ 
sr &ija.ija2015.homework2.game.HumanPlayer�҂��R�  xq ~       sq ~    w   q ~ q ~ 5xuq ~ :   q ~ %q ~ "q ~ sq ~ sq ~     w    x